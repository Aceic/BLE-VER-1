library verilog;
use verilog.vl_types.all;
entity dut is
end dut;
