package ovc_pkg;
	import ovm_pkg::*;
  import ovm_container_pkg::*;

`include "ovm_macros.svh"
`include "uvm_reg_macros.svh"
  import uvm_reg_pkg::*;
 import ble_reg_bank_pkg::*;

`include "tb_defs.sv"


`include "ahb_seq_item.sv"
 `include "ahb_coverage.sv"
//`include "adv_seq_item.sv"

`include "ahb_adapter.svh"
`include "ahb_agent_config.sv"
//`include "ahb_env_config.sv"
`include "ble_ovc_config.sv"
`include "ahb_master_driver.sv"
`include "ahb_master_monitor.sv"
`include "ahb_master_sequencer.sv"
`include "ahb_master_agent.sv"
//`include "ahb_scoreboard.sv"
//`include "ahb_master_uvc.sv"
//`include "ahb_seq.sv"
`include "ble_base_seq.sv"
`include "ble_ovc.sv"
`include "ble_ovc_virtual_seq.sv"



endpackage
