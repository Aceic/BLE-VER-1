library verilog;
use verilog.vl_types.all;
entity soc is
    port(
        rst             : in     vl_logic
    );
end soc;
