

interface intr_if();

 logic int_o;
 
endinterface
