`include "adv_config_test.sv"
