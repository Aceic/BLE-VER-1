`include "vip_define.sv"
// State register
`define status_register             `rstatus_register

// ADV state register 

`define adv_types                         `radv_types	                 	                   
`define adv_source_device_addr_lsb	      `radv_source_device_addr_lsb
`define adv_source_device_addr_msb	      `radv_source_device_addr_msb
`define adv_target_device_addr_lsb	      `radv_target_device_addr_lsb
`define adv_target_device_addr_msb	      `radv_target_device_addr_msb
`define adv_TX_Data	                      `radv_TX_Data	              
`define adv_RX_Data	                      `radv_RX_Data	              
`define adv_interval	                    `radv_interval	            
`define adv_interval_min	                `radv_interval_min	        
`define adv_interval_max	                `radv_interval_max	        
`define adv_channel_map_lsb	              `radv_channel_map_lsb	      
`define adv_channel_map_msb	              `radv_channel_map_msb	      
`define whitelist_reg	                    `rwhitelist_reg	            
`define adv_rx_type	                      `radv_rx_type	              


