

interface channel_if();

 
 logic [39:0] channel;

 
endinterface
