package vip_pkg;

   import ovm_pkg::*;
   import ovm_container_pkg::*;
   import uvm_reg_pkg::*;
   `include "uvm_reg_macros.svh"
   import ble_reg_bank_pkg::*;
   `include "ovm_macros.svh"

  // import tx_agent_pkg::*;
    import ahb_slv_pkg::*;
    import ctrl_pkg::*;
   

  

  `include "ble_vip_config.sv"
  `include "vip_env.sv"  
 





endpackage
